module top #(
    parameter CLK_F = 100_000_000
) (
    ports
);
    
endmodule