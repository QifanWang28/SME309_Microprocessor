module top_display_rom (
    input btn_p,
    input btn_spdup,
    input btn_spddn,
    input clk,
    output [7:0] anode,
    output [6:0] cathode,
    output dp,
    output [7:0] led
);
    
endmodule