module Cache (
    input [31:0] Addr,
    
    output hit,
    output [31:0] data
);
    
endmodule   